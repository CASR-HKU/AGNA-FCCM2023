`ifndef PARAM_SV
`define PARAM_SV

`define HW_DSP_CASCADED
`define HW_CONFIG_PE_NUM 21
`define HW_CONFIG_A_K 1
`define HW_CONFIG_A_C 8
`define HW_CONFIG_A_I 1
`define HW_CONFIG_A_J 1
`define HW_CONFIG_A_H 2
`define HW_CONFIG_A_W 13
`define HW_CONFIG_MACC_WIDTH 8

`endif
